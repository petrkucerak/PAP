module adder_full(
   input [31:0] a;
   input [31:0] b;
   output [31:0] c;
)
   // TODO: implement it
endmodule